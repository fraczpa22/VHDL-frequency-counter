-------------------------------------------------------------------------------
--
-- Title       : Fub1
-- Design      : TOP
-- Author      : IE
-- Company     : AGH
--
-------------------------------------------------------------------------------
--
-- File        : C:/My_Designs/TOP/TOP/src/Fub1.vhd
-- Generated   : Wed Jan 26 10:08:31 2022
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {Fub1} architecture {Fub1}}



entity Fub1 is
end Fub1;

--}} End of automatically maintained section

architecture Fub1 of Fub1 is
begin

	 -- enter your statements here --

end Fub1;
