library ieee;
use ieee.STD_LOGIC_UNSIGNED.all;
use ieee.std_logic_1164.all;

	-- Add your library and packages declaration here ...

entity kaskada_liczaca_TB is
end kaskada_liczaca_TB;

architecture TB_ARCHITECTURE of kaskada_liczaca_TB is
	-- Component declaration of the tested unit
	-- Component declaration of the tested unit
	component kaskada_liczaca
	port(
		CLK : in STD_LOGIC;
		CE : in STD_LOGIC;
		CLR : in STD_LOGIC;
		bit_wej : in STD_LOGIC;
		bity_wyj : out std_logic_vector(15 downto 0)
		);	
	end component;
	
		signal CLK : STD_LOGIC:= '0'; 
		signal CE : STD_LOGIC:= '0';
 		signal CLR: STD_LOGIC:= '1';
		signal bit_wej: STD_LOGIC:= '0'; 
		signal bity_wyj: STD_LOGIC_VECTOR(15 downto 0):=(others=>'0'); 
		signal bit_spr: STD_LOGIC_VECTOR(15 downto 0):=(others=>'0'); 
		--signal jaki_stan: STD_LOGIC_VECTOR(1 downto 0);

	constant period : time := 25 ns;

	-- Add your code here ...

begin

	-- Unit Under Test port map
	UUT : kaskada_liczaca
	port map (
			CLK=>CLK,
			CE=>CE,
			CLR => CLR,
			bit_wej => bit_wej,
 			bity_wyj => bity_wyj
			--jaki_stan=>jaki_stan
		);

CLOCK_CLK : process
begin
		CLK <= '0';
		wait for period/8; --0 fs
		CLK <= '1';
		wait for period/8; --50 ns
end process;

	
simul_1 : process
begin 
	CE<='1';
	CLR<='0';
	bit_wej<='0';	
	wait for period;
	bit_wej<='1';
	bit_spr<=bit_spr+1;
	wait for period; 
	bit_wej<='0';	
	wait for period;


end process; 




	-- Add your stimulus here ...

end TB_ARCHITECTURE;

configuration TESTBENCH_FOR_kaskada_liczaca of kaskada_liczaca_TB is
	for TB_ARCHITECTURE
		for UUT : kaskada_liczaca
			use entity work.kaskada_liczaca(kaskada_liczaca);
		end for;
	end for;
end TESTBENCH_FOR_kaskada_liczaca;

